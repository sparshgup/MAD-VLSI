magic
tech sky130A
timestamp 1759609458
<< nwell >>
rect -20 210 185 350
<< nmos >>
rect 50 0 65 100
<< pmos >>
rect 50 230 65 330
<< ndiff >>
rect 0 85 50 100
rect 0 15 15 85
rect 35 15 50 85
rect 0 0 50 15
rect 65 85 115 100
rect 65 15 80 85
rect 100 15 115 85
rect 65 0 115 15
<< pdiff >>
rect 0 315 50 330
rect 0 245 15 315
rect 35 245 50 315
rect 0 230 50 245
rect 65 315 115 330
rect 65 245 80 315
rect 100 245 115 315
rect 65 230 115 245
<< ndiffc >>
rect 15 15 35 85
rect 80 15 100 85
<< pdiffc >>
rect 15 245 35 315
rect 80 245 100 315
<< psubdiff >>
rect 115 85 165 100
rect 115 15 130 85
rect 150 15 165 85
rect 115 0 165 15
<< nsubdiff >>
rect 115 315 165 330
rect 115 245 130 315
rect 150 245 165 315
rect 115 230 165 245
<< psubdiffcont >>
rect 130 15 150 85
<< nsubdiffcont >>
rect 130 245 150 315
<< poly >>
rect 125 465 185 475
rect 125 445 135 465
rect 155 460 185 465
rect 155 445 165 460
rect 125 435 165 445
rect 50 330 65 345
rect 50 175 65 230
rect 50 165 90 175
rect 50 145 60 165
rect 80 145 90 165
rect 50 135 90 145
rect 50 100 65 135
rect 50 -15 65 0
rect 125 -85 165 -75
rect 125 -105 135 -85
rect 155 -100 165 -85
rect 155 -105 185 -100
rect 125 -115 185 -105
<< polycont >>
rect 135 445 155 465
rect 60 145 80 165
rect 135 -105 155 -85
<< locali >>
rect 125 465 165 475
rect 125 455 135 465
rect 25 445 135 455
rect 155 445 165 465
rect 25 435 165 445
rect 25 325 45 435
rect 5 315 45 325
rect 5 245 15 315
rect 35 245 45 315
rect 5 235 45 245
rect 70 315 160 325
rect 70 245 80 315
rect 100 245 130 315
rect 150 245 160 315
rect 70 235 160 245
rect 5 95 25 235
rect 50 165 90 175
rect 50 145 60 165
rect 80 155 90 165
rect 145 165 185 175
rect 145 155 155 165
rect 80 145 155 155
rect 175 145 185 165
rect 50 135 185 145
rect 5 85 45 95
rect 5 15 15 85
rect 35 15 45 85
rect 5 5 45 15
rect 70 85 160 95
rect 70 15 80 85
rect 100 15 130 85
rect 150 15 160 85
rect 70 5 160 15
rect 25 -75 45 5
rect 25 -85 165 -75
rect 25 -95 135 -85
rect 125 -105 135 -95
rect 155 -105 165 -85
rect 125 -115 165 -105
<< viali >>
rect 80 245 100 315
rect 130 245 150 315
rect 60 145 80 165
rect 155 145 175 165
rect 80 15 100 85
rect 130 15 150 85
<< metal1 >>
rect -20 315 185 586
rect -20 245 80 315
rect 100 245 130 315
rect 150 245 185 315
rect -20 230 185 245
rect -20 165 90 175
rect -20 145 60 165
rect 80 145 90 165
rect -20 135 90 145
rect 145 165 185 175
rect 145 145 155 165
rect 175 145 185 165
rect 145 135 185 145
rect -20 85 185 100
rect -20 15 80 85
rect 100 15 130 85
rect 150 15 185 85
rect -20 -246 185 15
rect -20 -340 185 -300
<< labels >>
rlabel metal1 81 582 81 582 1 VDD
rlabel metal1 82 -245 82 -245 1 GND
rlabel metal1 -19 154 -19 154 3 A
rlabel metal1 180 155 180 155 1 Y
<< end >>
