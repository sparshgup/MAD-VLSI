magic
tech sky130A
timestamp 1758238523
<< nwell >>
rect -100 480 340 620
<< nmos >>
rect 140 0 180 100
<< pmos >>
rect 140 500 180 600
<< ndiff >>
rect 0 80 140 100
rect 0 20 20 80
rect 60 20 140 80
rect 0 0 140 20
rect 180 80 320 100
rect 180 20 260 80
rect 300 20 320 80
rect 180 0 320 20
<< pdiff >>
rect 0 580 140 600
rect 0 520 20 580
rect 60 520 140 580
rect 0 500 140 520
rect 180 580 320 600
rect 180 520 260 580
rect 300 520 320 580
rect 180 500 320 520
<< ndiffc >>
rect 20 20 60 80
rect 260 20 300 80
<< pdiffc >>
rect 20 520 60 580
rect 260 520 300 580
<< psubdiff >>
rect -80 80 0 100
rect -80 20 -60 80
rect -20 20 0 80
rect -80 0 0 20
<< nsubdiff >>
rect -80 580 0 600
rect -80 520 -60 580
rect -20 520 0 580
rect -80 500 0 520
<< psubdiffcont >>
rect -60 20 -20 80
<< nsubdiffcont >>
rect -60 520 -20 580
<< poly >>
rect 140 600 180 640
rect 140 310 180 500
rect -100 300 180 310
rect -100 280 -90 300
rect -70 280 180 300
rect -100 270 180 280
rect 140 100 180 270
rect 140 -20 180 0
<< polycont >>
rect -90 280 -70 300
<< locali >>
rect -70 580 70 590
rect -70 520 -60 580
rect -20 520 20 580
rect 60 520 70 580
rect -70 510 70 520
rect 250 580 310 590
rect 250 520 260 580
rect 300 520 310 580
rect 250 510 310 520
rect -100 300 -60 310
rect -100 280 -90 300
rect -70 280 -60 300
rect -100 270 -60 280
rect -70 80 70 90
rect -70 20 -60 80
rect -20 20 20 80
rect 60 20 70 80
rect -70 10 70 20
rect 250 80 310 90
rect 250 20 260 80
rect 300 20 310 80
rect 250 10 310 20
<< viali >>
rect 20 520 60 580
rect 260 520 300 580
rect -90 280 -70 300
rect 20 20 60 80
rect 260 20 300 80
<< metal1 >>
rect 0 670 320 730
rect 10 580 70 670
rect 10 520 20 580
rect 60 520 70 580
rect 10 510 70 520
rect 250 580 310 590
rect 250 520 260 580
rect 300 520 310 580
rect 250 320 310 520
rect -140 300 -60 310
rect -140 280 -90 300
rect -70 280 -60 300
rect -140 270 -60 280
rect 250 260 370 320
rect 10 80 70 90
rect 10 20 20 80
rect 60 20 70 80
rect 10 -50 70 20
rect 250 80 310 260
rect 250 20 260 80
rect 300 20 310 80
rect 250 10 310 20
rect 0 -110 320 -50
<< labels >>
rlabel metal1 316 700 317 702 1 VDD
rlabel metal1 315 -79 316 -77 1 GND
rlabel metal1 366 291 367 291 1 Y
port 2 n
rlabel metal1 -120 290 -120 290 1 A
port 1 n
<< end >>
