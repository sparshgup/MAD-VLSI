magic
tech sky130A
timestamp 1759602863
<< nwell >>
rect -70 570 490 985
<< nmos >>
rect 0 370 15 470
rect 40 370 55 470
rect 105 370 120 470
rect 270 370 285 470
rect 335 370 350 470
rect 400 370 415 470
rect 0 125 15 225
rect 40 125 55 225
rect 105 125 120 225
rect 270 125 285 225
rect 335 125 350 225
rect 400 125 415 225
<< pmos >>
rect 0 855 15 955
rect 65 855 80 955
rect 130 855 145 955
rect 295 855 310 955
rect 335 855 350 955
rect 400 855 415 955
rect 0 600 15 700
rect 65 600 80 700
rect 130 600 145 700
rect 295 600 310 700
rect 335 600 350 700
rect 400 600 415 700
<< ndiff >>
rect -50 455 0 470
rect -50 385 -35 455
rect -15 385 0 455
rect -50 370 0 385
rect 15 370 40 470
rect 55 455 105 470
rect 55 385 70 455
rect 90 385 105 455
rect 55 370 105 385
rect 120 455 170 470
rect 120 385 135 455
rect 155 385 170 455
rect 120 370 170 385
rect 220 455 270 470
rect 220 385 235 455
rect 255 385 270 455
rect 220 370 270 385
rect 285 455 335 470
rect 285 385 300 455
rect 320 385 335 455
rect 285 370 335 385
rect 350 455 400 470
rect 350 385 365 455
rect 385 385 400 455
rect 350 370 400 385
rect 415 455 465 470
rect 415 385 430 455
rect 450 385 465 455
rect 415 370 465 385
rect -50 210 0 225
rect -50 140 -35 210
rect -15 140 0 210
rect -50 125 0 140
rect 15 125 40 225
rect 55 210 105 225
rect 55 140 70 210
rect 90 140 105 210
rect 55 125 105 140
rect 120 210 170 225
rect 120 140 135 210
rect 155 140 170 210
rect 120 125 170 140
rect 220 210 270 225
rect 220 140 235 210
rect 255 140 270 210
rect 220 125 270 140
rect 285 210 335 225
rect 285 140 300 210
rect 320 140 335 210
rect 285 125 335 140
rect 350 210 400 225
rect 350 140 365 210
rect 385 140 400 210
rect 350 125 400 140
rect 415 210 465 225
rect 415 140 430 210
rect 450 140 465 210
rect 415 125 465 140
<< pdiff >>
rect -50 940 0 955
rect -50 870 -35 940
rect -15 870 0 940
rect -50 855 0 870
rect 15 940 65 955
rect 15 870 30 940
rect 50 870 65 940
rect 15 855 65 870
rect 80 940 130 955
rect 80 870 95 940
rect 115 870 130 940
rect 80 855 130 870
rect 145 940 195 955
rect 145 870 160 940
rect 180 870 195 940
rect 145 855 195 870
rect 245 940 295 955
rect 245 870 260 940
rect 280 870 295 940
rect 245 855 295 870
rect 310 855 335 955
rect 350 940 400 955
rect 350 870 365 940
rect 385 870 400 940
rect 350 855 400 870
rect 415 940 465 955
rect 415 870 430 940
rect 450 870 465 940
rect 415 855 465 870
rect -50 685 0 700
rect -50 615 -35 685
rect -15 615 0 685
rect -50 600 0 615
rect 15 685 65 700
rect 15 615 30 685
rect 50 615 65 685
rect 15 600 65 615
rect 80 685 130 700
rect 80 615 95 685
rect 115 615 130 685
rect 80 600 130 615
rect 145 685 195 700
rect 145 615 160 685
rect 180 615 195 685
rect 145 600 195 615
rect 245 685 295 700
rect 245 615 260 685
rect 280 615 295 685
rect 245 600 295 615
rect 310 600 335 700
rect 350 685 400 700
rect 350 615 365 685
rect 385 615 400 685
rect 350 600 400 615
rect 415 685 465 700
rect 415 615 430 685
rect 450 615 465 685
rect 415 600 465 615
<< ndiffc >>
rect -35 385 -15 455
rect 70 385 90 455
rect 135 385 155 455
rect 235 385 255 455
rect 300 385 320 455
rect 365 385 385 455
rect 430 385 450 455
rect -35 140 -15 210
rect 70 140 90 210
rect 135 140 155 210
rect 235 140 255 210
rect 300 140 320 210
rect 365 140 385 210
rect 430 140 450 210
<< pdiffc >>
rect -35 870 -15 940
rect 30 870 50 940
rect 95 870 115 940
rect 160 870 180 940
rect 260 870 280 940
rect 365 870 385 940
rect 430 870 450 940
rect -35 615 -15 685
rect 30 615 50 685
rect 95 615 115 685
rect 160 615 180 685
rect 260 615 280 685
rect 365 615 385 685
rect 430 615 450 685
<< psubdiff >>
rect 220 320 320 335
rect 220 300 235 320
rect 305 300 320 320
rect 220 285 320 300
<< nsubdiff >>
rect -50 785 50 800
rect -50 765 -35 785
rect 35 765 50 785
rect -50 750 50 765
<< psubdiffcont >>
rect 235 300 305 320
<< nsubdiffcont >>
rect -35 765 35 785
<< poly >>
rect 375 1000 415 1010
rect 375 980 385 1000
rect 405 980 415 1000
rect 375 970 415 980
rect 0 955 15 970
rect 65 955 80 970
rect 130 955 145 970
rect 295 955 310 970
rect 335 955 350 970
rect 400 955 415 970
rect 0 840 15 855
rect -60 825 15 840
rect 0 700 15 715
rect 65 700 80 855
rect 130 840 145 855
rect 295 840 310 855
rect 105 830 145 840
rect 105 810 115 830
rect 135 810 145 830
rect 105 800 145 810
rect 170 830 310 840
rect 170 810 180 830
rect 200 825 310 830
rect 200 810 210 825
rect 170 800 210 810
rect 170 730 185 800
rect 130 715 185 730
rect 130 700 145 715
rect 295 700 310 715
rect 335 700 350 855
rect 400 840 415 855
rect 440 825 490 840
rect 440 755 455 825
rect 375 745 455 755
rect 375 725 385 745
rect 405 740 455 745
rect 405 725 415 740
rect 375 715 415 725
rect 400 700 415 715
rect 0 545 15 600
rect 65 585 80 600
rect 130 585 145 600
rect 295 585 310 600
rect -25 535 15 545
rect -25 515 -15 535
rect 5 515 15 535
rect -25 505 15 515
rect 0 470 15 505
rect 40 570 80 585
rect 105 570 145 585
rect 270 575 310 585
rect 40 470 55 570
rect 105 470 120 570
rect 270 555 280 575
rect 300 555 310 575
rect 270 545 310 555
rect 270 470 285 545
rect 335 470 350 600
rect 400 470 415 600
rect 0 355 15 370
rect -60 240 15 255
rect 0 225 15 240
rect 40 225 55 370
rect 105 355 120 370
rect 270 355 285 370
rect 80 344 120 355
rect 80 325 90 344
rect 110 330 120 344
rect 110 325 160 330
rect 80 315 160 325
rect 145 255 160 315
rect 145 240 285 255
rect 105 225 120 240
rect 270 225 285 240
rect 335 225 350 370
rect 400 355 415 370
rect 400 340 455 355
rect 440 280 455 340
rect 375 270 415 280
rect 375 250 385 270
rect 405 250 415 270
rect 375 240 415 250
rect 440 270 480 280
rect 440 250 450 270
rect 470 255 480 270
rect 470 250 490 255
rect 440 240 490 250
rect 400 225 415 240
rect 0 110 15 125
rect 40 70 55 125
rect 105 110 120 125
rect 270 110 285 125
rect 80 100 120 110
rect 80 80 90 100
rect 110 80 120 100
rect 80 70 120 80
rect 335 70 350 125
rect 400 110 415 125
rect 15 60 55 70
rect 15 40 25 60
rect 45 40 55 60
rect 15 30 55 40
rect 310 60 350 70
rect 310 40 320 60
rect 340 40 350 60
rect 310 30 350 40
<< polycont >>
rect 385 980 405 1000
rect 115 810 135 830
rect 180 810 200 830
rect 385 725 405 745
rect -15 515 5 535
rect 280 555 300 575
rect 90 325 110 344
rect 385 250 405 270
rect 450 250 470 270
rect 90 80 110 100
rect 25 40 45 60
rect 320 40 340 60
<< locali >>
rect 375 1000 415 1010
rect 375 990 385 1000
rect -24 970 104 990
rect -24 950 -5 970
rect 85 950 104 970
rect 315 980 385 990
rect 405 980 415 1000
rect 315 970 415 980
rect -45 940 -5 950
rect -45 870 -35 940
rect -15 870 -5 940
rect -45 860 -5 870
rect 20 940 60 950
rect 20 870 30 940
rect 50 870 60 940
rect 20 860 60 870
rect 85 940 125 950
rect 85 870 95 940
rect 115 870 125 940
rect 85 860 125 870
rect 150 940 190 950
rect 150 870 160 940
rect 180 870 190 940
rect 150 860 190 870
rect 20 795 40 860
rect 170 840 190 860
rect 250 940 290 950
rect 250 870 260 940
rect 280 870 290 940
rect 250 860 290 870
rect 105 830 145 840
rect 105 810 115 830
rect 135 810 145 830
rect 105 800 145 810
rect 170 830 210 840
rect 170 810 180 830
rect 200 810 210 830
rect 170 800 210 810
rect -45 785 45 795
rect -45 765 -35 785
rect 35 765 45 785
rect -45 755 45 765
rect 20 695 40 755
rect 125 750 145 800
rect 125 730 170 750
rect 150 695 170 730
rect 250 695 270 860
rect 315 695 335 970
rect 355 940 395 950
rect 355 870 365 940
rect 385 870 395 940
rect 355 860 395 870
rect 420 940 460 950
rect 420 870 430 940
rect 450 870 460 940
rect 420 860 460 870
rect 375 755 395 860
rect 375 745 415 755
rect 375 725 385 745
rect 405 725 415 745
rect 375 715 415 725
rect 440 695 460 860
rect -45 685 -5 695
rect -45 615 -35 685
rect -15 615 -5 685
rect -45 605 -5 615
rect 20 685 60 695
rect 20 615 30 685
rect 50 615 60 685
rect 20 605 60 615
rect 85 685 125 695
rect 85 615 95 685
rect 115 615 125 685
rect 85 605 125 615
rect 150 685 190 695
rect 150 615 160 685
rect 180 615 190 685
rect 150 605 190 615
rect 250 685 290 695
rect 250 615 260 685
rect 280 615 290 685
rect 315 685 395 695
rect 315 675 365 685
rect 250 605 290 615
rect 355 615 365 675
rect 385 615 395 685
rect 355 605 395 615
rect 420 685 460 695
rect 420 615 430 685
rect 450 615 460 685
rect 420 605 460 615
rect -25 585 -5 605
rect 85 585 105 605
rect -25 565 105 585
rect 150 585 170 605
rect 375 585 395 605
rect 150 575 310 585
rect 150 565 280 575
rect -25 535 15 545
rect -25 525 -15 535
rect -60 515 -15 525
rect 5 515 15 535
rect 150 525 170 565
rect 270 555 280 565
rect 300 555 310 575
rect 375 565 460 585
rect 270 545 310 555
rect -60 505 15 515
rect 80 505 170 525
rect 440 505 460 565
rect 80 465 100 505
rect 245 485 375 505
rect 245 465 265 485
rect 355 465 375 485
rect 440 485 490 505
rect 440 465 460 485
rect -45 455 -5 465
rect -45 385 -35 455
rect -15 385 -5 455
rect 60 455 100 465
rect 60 395 70 455
rect -45 375 -5 385
rect 20 385 70 395
rect 90 385 100 455
rect 20 375 100 385
rect 125 455 165 465
rect 125 385 135 455
rect 155 385 165 455
rect 125 375 165 385
rect 225 455 265 465
rect 225 385 235 455
rect 255 385 265 455
rect 225 375 265 385
rect 290 455 330 465
rect 290 385 300 455
rect 320 385 330 455
rect 290 375 330 385
rect 355 455 395 465
rect 355 385 365 455
rect 385 385 395 455
rect 355 375 395 385
rect 420 455 460 465
rect 420 385 430 455
rect 450 385 460 455
rect 420 375 460 385
rect -45 220 -25 375
rect -45 210 -5 220
rect -45 140 -35 210
rect -15 140 -5 210
rect -45 130 -5 140
rect 20 110 40 375
rect 80 344 120 355
rect 80 325 90 344
rect 110 325 120 344
rect 80 315 120 325
rect 80 220 100 315
rect 145 220 165 375
rect 290 330 310 375
rect 420 355 440 375
rect 395 335 440 355
rect 225 320 315 330
rect 225 300 235 320
rect 305 300 315 320
rect 225 290 315 300
rect 290 220 310 290
rect 395 280 415 335
rect 375 270 415 280
rect 375 250 385 270
rect 405 250 415 270
rect 375 240 415 250
rect 440 270 480 280
rect 440 250 450 270
rect 470 250 480 270
rect 440 240 480 250
rect 440 220 460 240
rect 60 210 100 220
rect 60 140 70 210
rect 90 140 100 210
rect 60 130 100 140
rect 125 210 165 220
rect 125 140 135 210
rect 155 140 165 210
rect 125 130 165 140
rect 225 210 265 220
rect 225 140 235 210
rect 255 140 265 210
rect 225 130 265 140
rect 290 210 330 220
rect 290 140 300 210
rect 320 140 330 210
rect 290 130 330 140
rect 355 210 395 220
rect 355 140 365 210
rect 385 140 395 210
rect 355 130 395 140
rect 420 210 460 220
rect 420 140 430 210
rect 450 140 460 210
rect 420 130 460 140
rect 245 110 265 130
rect 355 110 375 130
rect 20 100 120 110
rect 20 90 90 100
rect 80 80 90 90
rect 110 80 120 100
rect 245 90 375 110
rect 80 70 120 80
rect 15 60 55 70
rect 15 40 25 60
rect 45 40 55 60
rect 15 30 55 40
rect 310 60 350 70
rect 310 40 320 60
rect 340 40 350 60
rect 310 30 350 40
<< viali >>
rect 30 870 50 940
rect 260 870 280 940
rect -35 765 35 785
rect 430 870 450 940
rect 30 615 50 685
rect 260 615 280 685
rect 430 615 450 685
rect -35 385 -15 455
rect 135 385 155 455
rect 300 385 320 455
rect -35 140 -15 210
rect 235 300 305 320
rect 135 140 155 210
rect 300 140 320 210
rect 25 40 45 60
rect 320 40 340 60
<< metal1 >>
rect -60 940 490 956
rect -60 870 30 940
rect 50 870 260 940
rect 280 870 430 940
rect 450 870 490 940
rect -60 785 490 870
rect -60 765 -35 785
rect 35 765 490 785
rect -60 685 490 765
rect -60 615 30 685
rect 50 615 260 685
rect 280 615 430 685
rect 450 615 490 685
rect -60 600 490 615
rect -60 455 490 470
rect -60 385 -35 455
rect -15 385 135 455
rect 155 385 300 455
rect 320 385 490 455
rect -60 320 490 385
rect -60 300 235 320
rect 305 300 490 320
rect -60 210 490 300
rect -60 140 -35 210
rect -15 140 135 210
rect 155 140 300 210
rect 320 140 490 210
rect -60 124 490 140
rect -60 60 490 70
rect -60 40 25 60
rect 45 40 320 60
rect 340 40 490 60
rect -60 30 490 40
<< labels >>
rlabel metal1 -59 774 -59 774 7 VP
rlabel metal1 -59 307 -59 307 7 VN
rlabel metal1 -59 50 -59 50 7 CLK
rlabel locali -59 515 -59 515 7 D
rlabel poly -59 832 -59 832 7 Dn1
rlabel poly -59 247 -59 247 7 Dn2
rlabel locali 489 495 489 495 3 Q
rlabel poly 489 833 489 833 3 Qn
<< end >>
