magic
tech sky130A
timestamp 1759449554
<< nwell >>
rect -160 570 490 990
<< nmos >>
rect 0 260 15 360
rect 40 260 55 360
rect 105 260 120 360
rect 270 260 285 360
rect 335 260 350 360
rect 400 260 415 360
rect 0 0 15 100
rect 40 0 55 100
rect 105 0 120 100
rect 270 0 285 100
rect 335 0 350 100
rect 400 0 415 100
<< pmos >>
rect 0 860 15 960
rect 65 860 80 960
rect 130 860 145 960
rect 295 860 310 960
rect 335 860 350 960
rect 400 860 415 960
rect 0 600 15 700
rect 65 600 80 700
rect 130 600 145 700
rect 295 600 310 700
rect 335 600 350 700
rect 400 600 415 700
<< ndiff >>
rect -50 345 0 360
rect -50 275 -35 345
rect -15 275 0 345
rect -50 260 0 275
rect 15 260 40 360
rect 55 345 105 360
rect 55 275 70 345
rect 90 275 105 345
rect 55 260 105 275
rect 120 345 170 360
rect 120 275 135 345
rect 155 275 170 345
rect 120 260 170 275
rect 220 345 270 360
rect 220 275 235 345
rect 255 275 270 345
rect 220 260 270 275
rect 285 345 335 360
rect 285 275 300 345
rect 320 275 335 345
rect 285 260 335 275
rect 350 345 400 360
rect 350 275 365 345
rect 385 275 400 345
rect 350 260 400 275
rect 415 345 465 360
rect 415 275 430 345
rect 450 275 465 345
rect 415 260 465 275
rect -50 85 0 100
rect -50 15 -35 85
rect -15 15 0 85
rect -50 0 0 15
rect 15 0 40 100
rect 55 85 105 100
rect 55 15 70 85
rect 90 15 105 85
rect 55 0 105 15
rect 120 85 170 100
rect 120 15 135 85
rect 155 15 170 85
rect 120 0 170 15
rect 220 85 270 100
rect 220 15 235 85
rect 255 15 270 85
rect 220 0 270 15
rect 285 85 335 100
rect 285 15 300 85
rect 320 15 335 85
rect 285 0 335 15
rect 350 85 400 100
rect 350 15 365 85
rect 385 15 400 85
rect 350 0 400 15
rect 415 85 465 100
rect 415 15 430 85
rect 450 15 465 85
rect 415 0 465 15
<< pdiff >>
rect -50 945 0 960
rect -50 875 -35 945
rect -15 875 0 945
rect -50 860 0 875
rect 15 945 65 960
rect 15 875 30 945
rect 50 875 65 945
rect 15 860 65 875
rect 80 945 130 960
rect 80 875 95 945
rect 115 875 130 945
rect 80 860 130 875
rect 145 945 195 960
rect 145 875 160 945
rect 180 875 195 945
rect 145 860 195 875
rect 245 945 295 960
rect 245 875 260 945
rect 280 875 295 945
rect 245 860 295 875
rect 310 860 335 960
rect 350 945 400 960
rect 350 875 365 945
rect 385 875 400 945
rect 350 860 400 875
rect 415 945 465 960
rect 415 875 430 945
rect 450 875 465 945
rect 415 860 465 875
rect -50 685 0 700
rect -50 615 -35 685
rect -15 615 0 685
rect -50 600 0 615
rect 15 685 65 700
rect 15 615 30 685
rect 50 615 65 685
rect 15 600 65 615
rect 80 685 130 700
rect 80 615 95 685
rect 115 615 130 685
rect 80 600 130 615
rect 145 685 195 700
rect 145 615 160 685
rect 180 615 195 685
rect 145 600 195 615
rect 245 685 295 700
rect 245 615 260 685
rect 280 615 295 685
rect 245 600 295 615
rect 310 600 335 700
rect 350 685 400 700
rect 350 615 365 685
rect 385 615 400 685
rect 350 600 400 615
rect 415 685 465 700
rect 415 615 430 685
rect 450 615 465 685
rect 415 600 465 615
<< ndiffc >>
rect -35 275 -15 345
rect 70 275 90 345
rect 135 275 155 345
rect 235 275 255 345
rect 300 275 320 345
rect 365 275 385 345
rect 430 275 450 345
rect -35 15 -15 85
rect 70 15 90 85
rect 135 15 155 85
rect 235 15 255 85
rect 300 15 320 85
rect 365 15 385 85
rect 430 15 450 85
<< pdiffc >>
rect -35 875 -15 945
rect 30 875 50 945
rect 95 875 115 945
rect 160 875 180 945
rect 260 875 280 945
rect 365 875 385 945
rect 430 875 450 945
rect -35 615 -15 685
rect 30 615 50 685
rect 95 615 115 685
rect 160 615 180 685
rect 260 615 280 685
rect 365 615 385 685
rect 430 615 450 685
<< psubdiff >>
rect -140 85 -90 100
rect -140 15 -125 85
rect -105 15 -90 85
rect -140 0 -90 15
<< nsubdiff >>
rect -140 685 -90 700
rect -140 615 -125 685
rect -105 615 -90 685
rect -140 600 -90 615
<< psubdiffcont >>
rect -125 15 -105 85
<< nsubdiffcont >>
rect -125 615 -105 685
<< poly >>
rect 375 1005 415 1015
rect 375 985 385 1005
rect 405 985 415 1005
rect 375 975 415 985
rect 0 960 15 975
rect 65 960 80 975
rect 130 960 145 975
rect 295 960 310 975
rect 335 960 350 975
rect 400 960 415 975
rect 0 845 15 860
rect -50 830 15 845
rect 0 700 15 715
rect 65 700 80 860
rect 130 845 145 860
rect 295 845 310 860
rect 105 835 145 845
rect 105 815 115 835
rect 135 815 145 835
rect 105 805 145 815
rect 170 835 310 845
rect 170 815 180 835
rect 200 830 310 835
rect 200 815 210 830
rect 170 805 210 815
rect 170 730 185 805
rect 130 715 185 730
rect 130 700 145 715
rect 295 700 310 715
rect 335 700 350 860
rect 400 845 415 860
rect 440 830 490 845
rect 440 755 455 830
rect 375 745 455 755
rect 375 725 385 745
rect 405 740 455 745
rect 405 725 415 740
rect 375 715 415 725
rect 400 700 415 715
rect 0 450 15 600
rect 65 585 80 600
rect 130 585 145 600
rect 295 585 310 600
rect -25 440 15 450
rect -25 420 -15 440
rect 5 420 15 440
rect -25 410 15 420
rect 0 360 15 410
rect 40 570 80 585
rect 105 570 145 585
rect 270 575 310 585
rect 40 360 55 570
rect 105 360 120 570
rect 270 555 280 575
rect 300 555 310 575
rect 270 545 310 555
rect 270 360 285 545
rect 335 360 350 600
rect 400 360 415 600
rect 0 245 15 260
rect -50 115 15 130
rect 0 100 15 115
rect 40 100 55 260
rect 105 245 120 260
rect 270 245 285 260
rect 80 234 120 245
rect 80 215 90 234
rect 110 220 120 234
rect 110 215 160 220
rect 80 205 160 215
rect 145 130 160 205
rect 145 115 285 130
rect 105 100 120 115
rect 270 100 285 115
rect 335 100 350 260
rect 400 245 415 260
rect 400 230 455 245
rect 440 155 455 230
rect 375 145 415 155
rect 375 125 385 145
rect 405 125 415 145
rect 375 115 415 125
rect 440 145 480 155
rect 440 125 450 145
rect 470 130 480 145
rect 470 125 490 130
rect 440 115 490 125
rect 400 100 415 115
rect 0 -15 15 0
rect 40 -15 55 0
rect 105 -15 120 0
rect 270 -15 285 0
rect 335 -15 350 0
rect 400 -15 415 0
rect 80 -25 120 -15
rect 80 -45 90 -25
rect 110 -45 120 -25
rect 80 -55 120 -45
<< polycont >>
rect 385 985 405 1005
rect 115 815 135 835
rect 180 815 200 835
rect 385 725 405 745
rect -15 420 5 440
rect 280 555 300 575
rect 90 215 110 234
rect 385 125 405 145
rect 450 125 470 145
rect 90 -45 110 -25
<< locali >>
rect 375 1005 415 1015
rect 375 995 385 1005
rect -24 975 104 995
rect -24 955 -5 975
rect 85 955 104 975
rect 315 985 385 995
rect 405 985 415 1005
rect 315 975 415 985
rect -45 945 -5 955
rect -45 875 -35 945
rect -15 875 -5 945
rect -45 865 -5 875
rect 20 945 60 955
rect 20 875 30 945
rect 50 875 60 945
rect 20 865 60 875
rect 85 945 125 955
rect 85 875 95 945
rect 115 875 125 945
rect 85 865 125 875
rect 150 945 190 955
rect 150 875 160 945
rect 180 875 190 945
rect 150 865 190 875
rect 250 945 290 955
rect 250 875 260 945
rect 280 875 290 945
rect 250 865 290 875
rect 20 695 40 865
rect 170 845 190 865
rect 105 835 145 845
rect 105 815 115 835
rect 135 815 145 835
rect 105 805 145 815
rect 170 835 210 845
rect 170 815 180 835
rect 200 815 210 835
rect 170 805 210 815
rect 125 750 145 805
rect 125 730 170 750
rect 150 695 170 730
rect 315 695 335 975
rect 355 945 395 955
rect 355 875 365 945
rect 385 875 395 945
rect 355 865 395 875
rect 420 945 460 955
rect 420 875 430 945
rect 450 875 460 945
rect 420 865 460 875
rect 375 755 395 865
rect 375 745 415 755
rect 375 725 385 745
rect 405 725 415 745
rect 375 715 415 725
rect 440 695 460 865
rect -135 685 -95 695
rect -135 615 -125 685
rect -105 615 -95 685
rect -135 605 -95 615
rect -45 685 -5 695
rect -45 615 -35 685
rect -15 615 -5 685
rect -45 605 -5 615
rect 20 685 60 695
rect 20 615 30 685
rect 50 615 60 685
rect 20 605 60 615
rect 85 685 125 695
rect 85 615 95 685
rect 115 615 125 685
rect 85 605 125 615
rect 150 685 190 695
rect 150 615 160 685
rect 180 615 190 685
rect 150 605 190 615
rect 250 685 290 695
rect 250 615 260 685
rect 280 615 290 685
rect 315 685 395 695
rect 315 675 365 685
rect 250 605 290 615
rect 355 615 365 675
rect 385 615 395 685
rect 355 605 395 615
rect 420 685 460 695
rect 420 615 430 685
rect 450 615 460 685
rect 420 605 460 615
rect -25 585 -5 605
rect 85 585 105 605
rect -25 565 105 585
rect 150 585 170 605
rect 375 585 395 605
rect 150 575 310 585
rect 150 565 280 575
rect -25 440 15 450
rect -25 430 -15 440
rect -50 420 -15 430
rect 5 420 15 440
rect 150 430 170 565
rect 270 555 280 565
rect 300 555 310 575
rect 375 565 460 585
rect 270 545 310 555
rect -50 410 15 420
rect 80 410 170 430
rect 80 355 100 410
rect 440 395 460 565
rect 245 375 375 395
rect 245 355 265 375
rect 355 355 375 375
rect 440 375 490 395
rect 440 355 460 375
rect -45 345 -5 355
rect -45 275 -35 345
rect -15 275 -5 345
rect 60 345 100 355
rect 60 285 70 345
rect -45 265 -5 275
rect 20 275 70 285
rect 90 275 100 345
rect 20 265 100 275
rect 125 345 165 355
rect 125 275 135 345
rect 155 275 165 345
rect 125 265 165 275
rect 225 345 265 355
rect 225 275 235 345
rect 255 275 265 345
rect 225 265 265 275
rect 290 345 330 355
rect 290 275 300 345
rect 320 275 330 345
rect 290 265 330 275
rect 355 345 395 355
rect 355 275 365 345
rect 385 275 395 345
rect 355 265 395 275
rect 420 345 460 355
rect 420 275 430 345
rect 450 275 460 345
rect 420 265 460 275
rect -45 95 -25 265
rect -135 85 -95 95
rect -135 15 -125 85
rect -105 15 -95 85
rect -135 5 -95 15
rect -45 85 -5 95
rect -45 15 -35 85
rect -15 15 -5 85
rect -45 5 -5 15
rect 20 -15 40 265
rect 80 234 120 245
rect 80 215 90 234
rect 110 215 120 234
rect 80 205 120 215
rect 80 95 100 205
rect 145 95 165 265
rect 290 95 310 265
rect 420 245 440 265
rect 395 225 440 245
rect 395 155 415 225
rect 375 145 415 155
rect 375 125 385 145
rect 405 125 415 145
rect 375 115 415 125
rect 440 145 480 155
rect 440 125 450 145
rect 470 125 480 145
rect 440 115 480 125
rect 440 95 460 115
rect 60 85 100 95
rect 60 15 70 85
rect 90 15 100 85
rect 60 5 100 15
rect 125 85 165 95
rect 125 15 135 85
rect 155 15 165 85
rect 125 5 165 15
rect 225 85 265 95
rect 225 15 235 85
rect 255 15 265 85
rect 225 5 265 15
rect 290 85 330 95
rect 290 15 300 85
rect 320 15 330 85
rect 290 5 330 15
rect 355 85 395 95
rect 355 15 365 85
rect 385 15 395 85
rect 355 5 395 15
rect 420 85 460 95
rect 420 15 430 85
rect 450 15 460 85
rect 420 5 460 15
rect 245 -15 265 5
rect 355 -15 375 5
rect 20 -25 120 -15
rect 20 -35 90 -25
rect 80 -45 90 -35
rect 110 -45 120 -25
rect 245 -35 375 -15
rect 80 -55 120 -45
<< end >>
