magic
tech sky130A
timestamp 1758238574
<< nwell >>
rect -100 480 500 620
<< nmos >>
rect 100 0 140 100
rect 260 0 300 100
<< pmos >>
rect 100 500 140 600
rect 260 500 300 600
<< ndiff >>
rect 0 80 100 100
rect 0 20 20 80
rect 60 20 100 80
rect 0 0 100 20
rect 140 0 260 100
rect 300 80 400 100
rect 300 20 340 80
rect 380 20 400 80
rect 300 0 400 20
<< pdiff >>
rect 0 580 100 600
rect 0 520 20 580
rect 60 520 100 580
rect 0 500 100 520
rect 140 580 260 600
rect 140 520 180 580
rect 220 520 260 580
rect 140 500 260 520
rect 300 580 400 600
rect 300 520 340 580
rect 380 520 400 580
rect 300 500 400 520
<< ndiffc >>
rect 20 20 60 80
rect 340 20 380 80
<< pdiffc >>
rect 20 520 60 580
rect 180 520 220 580
rect 340 520 380 580
<< psubdiff >>
rect -80 80 0 100
rect -80 20 -60 80
rect -20 20 0 80
rect -80 0 0 20
<< nsubdiff >>
rect -80 580 0 600
rect -80 520 -60 580
rect -20 520 0 580
rect -80 500 0 520
rect 400 580 480 600
rect 400 520 420 580
rect 460 520 480 580
rect 400 500 480 520
<< psubdiffcont >>
rect -60 20 -20 80
<< nsubdiffcont >>
rect -60 520 -20 580
rect 420 520 460 580
<< poly >>
rect 100 600 140 640
rect 260 600 300 640
rect 100 410 140 500
rect 100 390 110 410
rect 130 390 140 410
rect 100 100 140 390
rect 260 200 300 500
rect 260 180 270 200
rect 290 180 300 200
rect 260 100 300 180
rect 100 -20 140 0
rect 260 -20 300 0
<< polycont >>
rect 110 390 130 410
rect 270 180 290 200
<< locali >>
rect -70 580 70 590
rect -70 520 -60 580
rect -20 520 20 580
rect 60 520 70 580
rect -70 510 70 520
rect 170 580 230 590
rect 170 520 180 580
rect 220 520 230 580
rect 170 510 230 520
rect 330 580 470 590
rect 330 520 340 580
rect 380 520 420 580
rect 460 520 470 580
rect 330 510 470 520
rect 100 410 140 420
rect 100 390 110 410
rect 130 390 140 410
rect 100 380 140 390
rect 260 200 300 210
rect 260 180 270 200
rect 290 180 300 200
rect 260 170 300 180
rect -70 80 70 90
rect -70 20 -60 80
rect -20 20 20 80
rect 60 20 70 80
rect -70 10 70 20
rect 330 80 390 90
rect 330 20 340 80
rect 380 20 390 80
rect 330 10 390 20
<< viali >>
rect 20 520 60 580
rect 180 520 220 580
rect 340 520 380 580
rect 110 390 130 410
rect 270 180 290 200
rect 20 20 60 80
rect 340 20 380 80
<< metal1 >>
rect 0 670 400 730
rect 10 580 70 670
rect 10 520 20 580
rect 60 520 70 580
rect 10 510 70 520
rect 170 580 230 590
rect 170 520 180 580
rect 220 520 230 580
rect -100 410 140 420
rect -100 390 110 410
rect 130 390 140 410
rect -100 380 140 390
rect 170 330 230 520
rect 330 580 390 670
rect 330 520 340 580
rect 380 520 390 580
rect 330 510 390 520
rect 170 260 500 330
rect -100 200 300 210
rect -100 180 270 200
rect 290 180 300 200
rect -100 170 300 180
rect 10 80 70 90
rect 10 20 20 80
rect 60 20 70 80
rect 10 -50 70 20
rect 330 80 390 260
rect 330 20 340 80
rect 380 20 390 80
rect 330 10 390 20
rect 0 -110 400 -50
<< labels >>
rlabel metal1 1 700 1 703 1 VDD
rlabel metal1 3 -84 3 -81 1 GND
rlabel metal1 -90 399 -89 400 1 A
port 2 n
rlabel metal1 -91 190 -90 191 1 B
port 1 n
rlabel metal1 360 299 361 300 1 Y
port 3 n
<< end >>
